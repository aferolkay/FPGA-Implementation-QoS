library verilog;
use verilog.vl_types.all;
entity deneme3_tb is
end deneme3_tb;
