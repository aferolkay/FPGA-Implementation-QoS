library verilog;
use verilog.vl_types.all;
entity deneme_tb is
end deneme_tb;
