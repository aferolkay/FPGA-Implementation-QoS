library verilog;
use verilog.vl_types.all;
entity deneme2_tb is
end deneme2_tb;
