library verilog;
use verilog.vl_types.all;
entity deneme4_tb is
end deneme4_tb;
